`timescale 1ns/1ns
module Shifters( A, S, R );

    input  [31:0] A;
    input  [4:0]  S;
    output [31:0] R;

endmodule
